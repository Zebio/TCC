module (
	input 
	output );

	wire hysteresis;
	assign hysteresis = ;


endmodule 
